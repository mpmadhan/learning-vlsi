//4:1 Decoder
//S0,S1 => selector bits
//D0,D1,D2,D3 => output values
module decoder(
  input S0,S1,D0,D1,D2,D3,
  output Y);

  assign Y = ; //decoder logic

endmodule    
